library verilog;
use verilog.vl_types.all;
entity control_test_vlg_vec_tst is
end control_test_vlg_vec_tst;
