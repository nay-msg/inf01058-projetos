library verilog;
use verilog.vl_types.all;
entity decod_vlg_vec_tst is
end decod_vlg_vec_tst;
