library verilog;
use verilog.vl_types.all;
entity mux8bits21_vlg_vec_tst is
end mux8bits21_vlg_vec_tst;
